package pkg;
	parameter MEM_DEPTH=512;
parameter ADDER_SIZE=8;
endpackage : pkg